* File: 3r3w.pex.netlist
* Created: Wed Sep 16 20:56:54 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt bitcell_3r3w  
+ W1_WL W2_WL W3_WL
+ ML1 ML2 ML3
+ W1_BTL W1_BTLB W2_BTL W2_BTLB W3_BTL W3_BTLB 
+ SL_1 SLB_1 SL_2 SLB_2 SL_3 SLB_3 
* 
MM0 GND! D Dbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 D Dbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM3 VDD! D Dbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 D Dbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM43 Dbar W3_WL W3_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM42 Dbar W2_WL W2_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM38 W3_BTL W3_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM39 W2_BTL W2_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM41 Dbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM40 W1_BTL W1_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM158 net0116 SL_2 GND! GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14
+ AS=2.835e-14 PD=8.2e-07 PS=7.5e-07
MM159 ML2 Dbar net0116 GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=3.78e-14
+ PD=7.5e-07 PS=8.2e-07
MM161 net0117 SL_3 GND! GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14
+ AS=2.835e-14 PD=8.2e-07 PS=7.5e-07
MM162 ML3 Dbar net0117 GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=3.78e-14
+ PD=7.5e-07 PS=8.2e-07
MM96 net109 SL_1 GND! GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
MM160 ML1 Dbar net109 GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=3.78e-14
+ PD=7.5e-07 PS=8.2e-07
MM167 net0177 SLB_3 GND! GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14
+ AS=2.835e-14 PD=8.2e-07 PS=7.5e-07
MM166 ML3 D net0177 GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=3.78e-14
+ PD=7.5e-07 PS=8.2e-07
MM171 net0179 SLB_1 GND! GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14
+ AS=2.835e-14 PD=8.2e-07 PS=7.5e-07
MM170 ML1 D net0179 GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=3.78e-14
+ PD=7.5e-07 PS=8.2e-07
MM168 net0172 SLB_2 GND! GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14
+ AS=2.835e-14 PD=8.2e-07 PS=7.5e-07
MM169 ML2 D net0172 GND! NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=3.78e-14
+ PD=7.5e-07 PS=8.2e-07
c_11 W1_BTLB 0 0.0570715f
c_22 W2_BTLB 0 0.0180055f
c_36 W3_BTLB 0 0.0240391f
c_54 W1_WL 0 0.0942915f
c_75 W3_WL 0 0.0868623f
c_95 W2_WL 0 0.0931474f
c_112 Dbar 0 0.26099f
c_126 SL_1 0 0.0644094f
c_143 SL_3 0 0.0876297f
c_157 SL_2 0 0.0645704f
c_175 ML1 0 0.0671055f
c_192 SLB_3 0 0.0910414f
c_206 SLB_2 0 0.064686f
c_223 D 0 0.261405f
c_237 SLB_1 0 0.0644094f
c_251 W3_BTL 0 0.0240848f
c_262 W1_BTL 0 0.0570715f
c_273 W2_BTL 0 0.0180055f
c_292 ML3 0 0.0456259f
c_312 ML2 0 0.0537474f
c_322 VDD! 0 0.0129674f
c_344 GND! 0 0.194289f
*
.include "3r3w.pex.netlist.3R3W.pxi"
*
.ends
*
*
