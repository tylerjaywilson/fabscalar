* File: 8r8w.pex.netlist
* Created: Sat Sep 12 11:30:35 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt bitcell_8r8w  
+ W1_WL W2_WL W3_WL W4_WL W5_WL W6_WL W7_WL W8_WL
+ ML1 ML2 ML3 ML4 ML5 ML6 ML7 ML8 
+ W1_BTL W1_BTLB W2_BTL W2_BTLB W3_BTL W3_BTLB W4_BTL W4_BTLB 
+ W5_BTL W5_BTLB W6_BTL W6_BTLB W7_BTL W7_BTLB W8_BTL W8_BTLB 
+ SL_1 SLB_1 SL_2 SLB_2 SL_3 SLB_3 SL_4 SLB_4 
+ SL_5 SLB_5 SL_6 SLB_6 SL_7 SLB_7 SL_8 SLB_8 
* 
MM3 VDD! D Dbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 D Dbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM43 Dbar W3_WL W3_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM55 Dbar W5_WL W5_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM41 Dbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM62 Dbar W7_WL W7_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM42 Dbar W2_WL W2_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM53 Dbar W4_WL W4_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM58 Dbar W6_WL W6_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM66 Dbar W8_WL W8_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM0 GND! D Dbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 D Dbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM59 W6_BTL W6_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM67 W8_BTL W8_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM38 W3_BTL W3_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM54 W5_BTL W5_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM40 W1_BTL W1_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM63 W7_BTL W7_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM39 W2_BTL W2_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM52 W4_BTL W4_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM128 net0116 SL_2 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM129 ML2 Dbar net0116 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM154 net0172 SLB_2 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM155 ML2 D net0172 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM136 net0131 SL_6 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM137 ML6 Dbar net0131 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM157 net0179 SLB_1 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM156 ML1 D net0179 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM153 net0177 SLB_3 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM152 ML3 D net0177 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM146 net0163 SLB_6 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM147 ML6 D net0163 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM150 net0128 SLB_4 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM151 ML4 D net0128 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM145 net0160 SLB_7 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM144 ML7 D net0160 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM149 net0167 SLB_5 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM148 ML5 D net0167 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM142 net0149 SLB_8 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM143 ML8 D net0149 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM96 net109 SL_1 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM127 ML1 Dbar net109 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM130 net0117 SL_3 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM131 ML3 Dbar net0117 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM133 net0124 SL_4 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM132 ML4 Dbar net0124 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM139 net0130 SL_7 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM138 ML7 Dbar net0130 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM135 net098 SL_5 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM134 ML5 Dbar net098 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM140 net0107 SL_8 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM141 ML8 Dbar net0107 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
c_25 W3_BTLB 0 0.0264926f
c_46 W1_BTLB 0 0.074191f
c_68 W2_BTLB 0 0.0328378f
c_108 W3_WL 0 0.11364f
c_151 W1_WL 0 0.106686f
c_192 W2_WL 0 0.105343f
c_233 W5_WL 0 0.0940433f
c_276 W7_WL 0 0.0983576f
c_317 W4_WL 0 0.100438f
c_344 W7_BTLB 0 0.0309722f
c_370 W4_BTLB 0 0.0331629f
c_396 W5_BTLB 0 0.0254827f
c_437 W6_WL 0 0.100939f
c_463 W6_BTLB 0 0.0250695f
c_492 SL_1 0 0.0735698f
c_522 SL_2 0 0.0740961f
c_561 Dbar 0 0.702987f
c_585 W8_BTLB 0 0.0197212f
c_612 SL_5 0 0.0722499f
c_636 SL_3 0 0.0743199f
c_662 SL_4 0 0.0647433f
c_686 SL_6 0 0.0689124f
c_711 SL_7 0 0.0784658f
c_752 ML6 0 0.0853511f
c_794 ML7 0 0.101033f
c_836 ML8 0 0.109155f
c_863 SL_8 0 0.128963f
c_890 SLB_8 0 0.129974f
c_915 SLB_7 0 0.0785111f
c_953 D 0 0.701611f
c_979 SLB_6 0 0.0689606f
c_1005 SLB_4 0 0.0647433f
c_1029 SLB_3 0 0.07432f
c_1056 SLB_5 0 0.0722645f
c_1080 W8_BTL 0 0.0197212f
c_1110 SLB_2 0 0.0740961f
c_1139 SLB_1 0 0.0735698f
c_1165 W6_BTL 0 0.0250695f
c_1191 W5_BTL 0 0.0254827f
c_1218 W7_BTL 0 0.0309722f
c_1244 W4_BTL 0 0.0331629f
c_1269 W3_BTL 0 0.0264926f
c_1290 W1_BTL 0 0.0736699f
c_1312 W2_BTL 0 0.0328378f
c_1353 W8_WL 0 0.108147f
c_1394 ML1 0 0.0620246f
c_1437 ML2 0 0.0666807f
c_1479 ML3 0 0.0649312f
c_1520 ML4 0 0.0697365f
c_1561 ML5 0 0.0750364f
c_1572 VDD! 0 0.0163964f
c_1626 GND! 0 0.693479f
c_1637 net0116 0 0.00897647f
c_1648 net0172 0 0.00897647f
*
.include "8r8w.pex.netlist.8R8W.pxi"
*
.ends
*
*
