* File: 8r4w_new.pex.netlist
* Created: Sun Oct 25 19:39:57 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
* 
.subckt bitcell_8r4w  R1_WL R2_WL R3_WL R4_WL R5_WL R6_WL R7_WL R8_WL
+ W1_WL W2_WL W3_WL W4_WL
+ R1_BTL R1_BTLB R2_BTL R2_BTLB R3_BTL R3_BTLB R4_BTL R4_BTLB
+ R5_BTL R5_BTLB R6_BTL R6_BTLB R7_BTL R7_BTLB R8_BTL R8_BTLB
+ W1_BTL W1_BTLB W2_BTL W2_BTLB W3_BTL W3_BTLB W4_BTL W4_BTLB

MM94 GND! qbar qbar_new GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM95 GND! q q_new GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM3 VDD! q qbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 q qbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM41 qbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM42 qbar W2_WL W2_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM43 qbar W3_WL W3_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM53 qbar W4_WL W4_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM47 R1_BTLB R1_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
MM48 R2_BTLB R2_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
MM40 W1_BTL W1_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM84 R7_BTL R7_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM85 R8_BTL R8_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM52 W4_BTL W4_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM39 W2_BTL W2_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM38 W3_BTL W3_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM49 R3_BTLB R3_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM60 R6_BTLB R6_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM51 R4_BTLB R4_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM65 R7_BTLB R7_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM57 R5_BTLB R5_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM68 R8_BTLB R8_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM0 GND! q qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 q qbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM81 R3_BTL R3_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM82 R6_BTL R6_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM78 R1_BTL R1_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM80 R4_BTL R4_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM79 R2_BTL R2_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM83 R5_BTL R5_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
c_19 W1_BTLB 0 0.0562849f
c_37 W2_BTLB 0 0.0212375f
c_57 W3_BTLB 0 0.0183189f
c_94 W1_WL 0 0.120703f
c_134 W2_WL 0 0.118176f
c_166 W3_WL 0 0.156049f
c_201 W4_WL 0 0.102496f
c_237 R1_WL 0 0.0969325f
c_272 R2_WL 0 0.104305f
c_292 R1_BTLB 0 0.0226724f
c_314 W4_BTLB 0 0.0294309f
c_335 R2_BTLB 0 0.0231715f
c_356 R3_BTLB 0 0.0234137f
c_376 R4_BTLB 0 0.0248016f
c_399 R5_BTLB 0 0.0240057f
c_433 R3_WL 0 0.0891297f
c_469 R4_WL 0 0.0838564f
c_503 R5_WL 0 0.0887066f
c_537 R6_WL 0 0.088602f
c_572 R7_WL 0 0.0778897f
c_607 R8_WL 0 0.0801927f
c_628 R6_BTLB 0 0.0240885f
c_650 R7_BTLB 0 0.0211531f
c_673 R8_BTLB 0 0.0234056f
c_694 R3_BTL 0 0.0220462f
c_717 R1_BTL 0 0.0232274f
c_739 R2_BTL 0 0.0210921f
c_760 R6_BTL 0 0.0240189f
c_782 R4_BTL 0 0.023751f
c_803 R5_BTL 0 0.0234729f
c_824 R7_BTL 0 0.022209f
c_844 R8_BTL 0 0.0214949f
c_866 W1_BTL 0 0.0292541f
c_885 W4_BTL 0 0.0230875f
c_905 W2_BTL 0 0.0183717f
c_923 W3_BTL 0 0.0563437f
c_948 qbar_new 0 0.0940928f
c_977 qbar 0 0.198031f
c_1015 GND! 0 0.16388f
c_1048 VDD! 0 0.134597f
c_1073 q_new 0 0.093468f
c_1102 q 0 0.193268f
*
.include "8r4w_new.pex.netlist.8R4W_NEW.pxi"
*
.ends
*
*
