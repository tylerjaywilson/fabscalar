* File: 1r1w.pex.netlist
* Created: Wed Sep 16 20:59:15 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt bitcell_1r1w  
+ W1_WL ML1
+ W1_BTL W1_BTLB SL_1 SLB_1
* 
MM0 GND! D Dbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 D Dbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM3 VDD! D Dbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 D Dbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM41 Dbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM40 W1_BTL W1_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM96 net109 SL_1 GND! GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM160 ML1 Dbar net109 GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM170 ML1 D net0179 GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM171 net0179 SLB_1 GND! GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
c_6 W1_BTLB 0 0.0312435f
c_14 SL_1 0 0.0677325f
c_23 W1_WL 0 0.11647f
c_31 SLB_1 0 0.0677325f
c_38 W1_BTL 0 0.0312161f
c_47 Dbar 0 0.11137f
c_56 VDD! 0 0.020124f
c_65 D 0 0.104626f
c_75 GND! 0 0.103739f
c_84 ML1 0 0.0563103f
*
.include "1r1w.pex.netlist.1R1W.pxi"
*
.ends
*
*
