* File: 8r8w.pex.netlist
* Created: Sun Nov  1 18:22:24 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt bitcell_8r8w  R1_WL R2_WL R3_WL R4_WL R5_WL R6_WL R7_WL R8_WL W1_WL W2_WL W3_WL W4_WL W5_WL
+ W6_WL W7_WL  W8_WL R1_BTL R1_BTLB R2_BTL R2_BTLB R3_BTL R3_BTLB R4_BTL R4_BTLB
+ R5_BTL R5_BTLB R6_BTL R6_BTLB R7_BTL R7_BTLB R8_BTL R8_BTLB W1_BTL W1_BTLB
+ W2_BTL W2_BTLB W3_BTL W3_BTLB W4_BTL W4_BTLB W5_BTL W5_BTLB
+ W6_BTL W6_BTLB W7_BTL  W7_BTLB W8_BTL  W8_BTLB 
* 
MM96 qbar_new qbar GND! GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM94 GND! q q_new GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM3 VDD! q qbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 q qbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM0 GND! q qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 q qbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM41 qbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM55 qbar W5_WL W5_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM47 R1_BTLB R1_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM57 R5_BTLB R5_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM42 qbar W2_WL W2_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM58 qbar W6_WL W6_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM48 R2_BTLB R2_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM60 R6_BTLB R6_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM43 qbar W3_WL W3_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM62 qbar W7_WL W7_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM49 R3_BTLB R3_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM65 R7_BTLB R7_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM53 qbar W4_WL W4_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM66 qbar W8_WL W8_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM51 R4_BTLB R4_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM68 R8_BTLB R8_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM78 R1_BTL R1_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM83 R5_BTL R5_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM40 W1_BTL W1_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM54 W5_BTL W5_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM79 R2_BTL R2_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM82 R6_BTL R6_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM39 W2_BTL W2_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM59 W6_BTL W6_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM81 R3_BTL R3_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM84 R7_BTL R7_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM38 W3_BTL W3_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM63 W7_BTL W7_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM80 R4_BTL R4_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM85 R8_BTL R8_WL q_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM52 W4_BTL W4_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM67 W8_BTL W8_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
c_24 W1_BTLB 0 0.0765253f
c_49 W2_BTLB 0 0.0357215f
c_73 W3_BTLB 0 0.0338723f
c_97 W4_BTLB 0 0.0285148f
c_142 W1_WL 0 0.131243f
c_185 W2_WL 0 0.111163f
c_232 W3_WL 0 0.12786f
c_272 W4_WL 0 0.114814f
c_314 W5_WL 0 0.110149f
c_361 W6_WL 0 0.128459f
c_403 W7_WL 0 0.109422f
c_444 W8_WL 0 0.17158f
c_469 W6_BTLB 0 0.031896f
c_497 W5_BTLB 0 0.0232344f
c_522 W7_BTLB 0 0.0274946f
c_547 W8_BTLB 0 0.0354735f
c_575 R1_BTLB 0 0.0361047f
c_601 R2_BTLB 0 0.0343487f
c_626 R3_BTLB 0 0.0290521f
c_652 R4_BTLB 0 0.0289385f
c_694 R1_WL 0 0.108407f
c_738 R2_WL 0 0.0959377f
c_781 R3_WL 0 0.103501f
c_824 R4_WL 0 0.104564f
c_866 R5_WL 0 0.0996474f
c_910 R6_WL 0 0.101187f
c_954 R7_WL 0 0.0892775f
c_997 R8_WL 0 0.0908987f
c_1023 R5_BTLB 0 0.0293083f
c_1047 R6_BTLB 0 0.0271234f
c_1073 R7_BTLB 0 0.023117f
c_1100 R8_BTLB 0 0.0299726f
c_1128 R1_BTL 0 0.0340017f
c_1153 R3_BTL 0 0.0271561f
c_1179 R4_BTL 0 0.0286235f
c_1203 R2_BTL 0 0.0246351f
c_1227 R6_BTL 0 0.0290508f
c_1253 R5_BTL 0 0.0301903f
c_1279 R7_BTL 0 0.0331961f
c_1307 R8_BTL 0 0.0349626f
c_1333 W2_BTL 0 0.0265003f
c_1359 W3_BTL 0 0.0323178f
c_1387 W4_BTL 0 0.0197287f
c_1414 W1_BTL 0 0.0374153f
c_1440 W5_BTL 0 0.0271968f
c_1465 W6_BTL 0 0.033503f
c_1489 W8_BTL 0 0.0720644f
c_1514 W7_BTL 0 0.034183f
c_1540 qbar_new 0 0.0873459f
c_1579 qbar 0 0.22629f
c_1625 GND! 0 0.230928f
c_1665 VDD! 0 0.186768f
c_1691 q_new 0 0.0916346f
c_1728 q 0 0.217502f
*
.include "8r8w.pex.netlist.8R8W.pxi"
*
.ends
*
*
