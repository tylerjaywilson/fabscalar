* File: 2r2w.pex.netlist
* Created: Wed Sep 16 20:57:48 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt bitcell_2r2w  
+ W1_WL W2_WL ML1 ML2
+ W1_BTL W1_BTLB W2_BTL W2_BTLB
+ SL_1 SLB_1 SL_2 SLB_2
* 
MM0 GND! D Dbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 D Dbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM3 VDD! D Dbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 D Dbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM158 net0116 SL_2 GND! GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM159 ML2 Dbar net0116 GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM96 net109 SL_1 GND! GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM160 ML1 Dbar net109 GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM170 ML1 D net0179 GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM171 net0179 SLB_1 GND! GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
MM169 ML2 D net0172 GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM168 net0172 SLB_2 GND! GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
MM41 Dbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM42 Dbar W2_WL W2_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM39 W2_BTL W2_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM40 W1_BTL W1_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
c_10 W1_BTLB 0 0.0307017f
c_23 W1_WL 0 0.100689f
c_33 SL_1 0 0.0527595f
c_47 W2_WL 0 0.0719307f
c_60 SL_2 0 0.0563686f
c_70 W2_BTLB 0 0.0205522f
c_80 W2_BTL 0 0.0205527f
c_93 SLB_2 0 0.0556239f
c_103 SLB_1 0 0.0527475f
c_113 W1_BTL 0 0.0313288f
c_126 Dbar 0 0.160479f
c_134 VDD! 0 0.0133917f
c_147 D 0 0.162028f
c_163 GND! 0 0.148839f
c_176 ML2 0 0.0418353f
c_188 ML1 0 0.0512062f
*
.include "2r2w.pex.netlist.2R2W.pxi"
*
.ends
*
*
