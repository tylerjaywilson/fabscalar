* File: 5r5w.pex.netlist
* Created: Wed Sep 16 20:52:54 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt bitcell_5r5w  
+ W1_WL W2_WL W3_WL W4_WL W5_WL
+ ML1 ML2 ML3 ML4 ML5
+ W1_BTL W1_BTLB W2_BTL W2_BTLB W3_BTL W3_BTLB W4_BTL W4_BTLB 
+ W5_BTL W5_BTLB
+ SL_1 SLB_1 SL_2 SLB_2 SL_3 SLB_3 SL_4 SLB_4 
+ SL_5 SLB_5 
* 
MM3 VDD! D Dbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 D Dbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM96 net109 SL_1 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM127 ML1 Dbar net109 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM128 net0116 SL_2 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM129 ML2 Dbar net0116 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM133 net0124 SL_4 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM132 ML4 Dbar net0124 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM130 net0117 SL_3 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM131 ML3 Dbar net0117 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM135 net098 SL_5 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
MM134 ML5 Dbar net098 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM153 net0177 SLB_3 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM152 ML3 D net0177 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM149 net0167 SLB_5 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM148 ML5 D net0167 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM150 net0128 SLB_4 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM151 ML4 D net0128 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM157 net0179 SLB_1 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM156 ML1 D net0179 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM154 net0172 SLB_2 GND! GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14
+ AS=3.78e-14 PD=1e-06 PS=9.3e-07
MM155 ML2 D net0172 GND! NMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
MM42 Dbar W2_WL W2_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM53 Dbar W4_WL W4_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM41 Dbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM52 W4_BTL W4_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM39 W2_BTL W2_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM40 W1_BTL W1_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM43 Dbar W3_WL W3_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM55 Dbar W5_WL W5_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM0 GND! D Dbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 D Dbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM38 W3_BTL W3_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM54 W5_BTL W5_WL D GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
c_16 W2_BTLB 0 0.0210671f
c_46 W2_WL 0 0.0948536f
c_62 W1_BTLB 0 0.0644773f
c_81 W4_BTLB 0 0.0220635f
c_108 W4_WL 0 0.0991515f
c_138 W1_WL 0 0.0988888f
c_157 W3_BTLB 0 0.0249117f
c_184 W3_WL 0 0.0868027f
c_204 SL_2 0 0.0573546f
c_223 SL_1 0 0.0626449f
c_249 Dbar 0 0.422146f
c_267 W5_BTLB 0 0.0303878f
c_284 SL_3 0 0.0616409f
c_302 SL_4 0 0.0649929f
c_332 ML4 0 0.077933f
c_360 ML5 0 0.090482f
c_382 SL_5 0 0.108468f
c_404 SLB_5 0 0.112915f
c_422 SLB_4 0 0.0650914f
c_447 D 0 0.419013f
c_466 SLB_3 0 0.0625315f
c_484 W5_BTL 0 0.0303575f
c_503 SLB_1 0 0.0626679f
c_523 SLB_2 0 0.0573714f
c_542 W3_BTL 0 0.0249117f
c_561 W4_BTL 0 0.0220539f
c_577 W1_BTL 0 0.0643986f
c_593 W2_BTL 0 0.020747f
c_620 W5_WL 0 0.0922927f
c_649 ML3 0 0.0619123f
c_661 VDD! 0 0.0117337f
c_695 GND! 0 0.419345f
c_722 ML1 0 0.0426195f
c_750 ML2 0 0.047482f
*
.include "5r5w.pex.netlist.5R5W.pxi"
*
.ends
*
*
