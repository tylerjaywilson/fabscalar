* File: 5r5w.pex.netlist
* Created: Sun Nov  1 18:37:37 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt  bitcell_5r5w  R1_WL R2_WL R3_WL R4_WL R5_WL
+ W1_WL W2_WL W3_WL W4_WL W5_WL
+ R1_BTL R1_BTLB R2_BTL R2_BTLB R3_BTL R3_BTLB R4_BTL R4_BTLB R5_BTL R5_BTLB
+ W1_BTL W1_BTLB W2_BTL W2_BTLB W3_BTL W3_BTLB W4_BTL W4_BTLB W5_BTL W5_BTLB
* 
MM97 GND! qbar qbar_new GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM96 GND! q qnew GND! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM3 VDD! q qbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 q qbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM94 qbar W5_WL W5_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM49 R3_BTLB R3_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
MM81 R3_BTL R3_WL qnew GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM95 W5_BTL W5_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM0 GND! q qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 q qbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM41 qbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM43 qbar W3_WL W3_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM48 R2_BTLB R2_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM57 R5_BTLB R5_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM42 qbar W2_WL W2_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM60 W4_BTLB W4_WL qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM47 R1_BTLB R1_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM51 R4_BTLB R4_WL qbar_new GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15
+ AS=1.26e-14 PD=3.9e-07 PS=4.6e-07
MM79 R2_BTL R2_WL qnew GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM83 R5_BTL R5_WL qnew GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM38 W3_BTL W3_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM40 W1_BTL W1_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM78 R1_BTL R1_WL qnew GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM80 R4_BTL R4_WL qnew GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM82 W4_BTL W4_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM39 W2_BTL W2_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
c_16 W1_BTLB 0 0.047076f
c_33 W2_BTLB 0 0.0247044f
c_66 W1_WL 0 0.10851f
c_98 W2_WL 0 0.110493f
c_128 W3_WL 0 0.0860364f
c_158 W4_WL 0 0.090598f
c_184 W5_WL 0 0.131827f
c_203 W4_BTLB 0 0.0209705f
c_222 W3_BTLB 0 0.0228965f
c_241 W5_BTLB 0 0.0257566f
c_262 R2_BTLB 0 0.0233371f
c_281 R1_BTLB 0 0.0230702f
c_311 R2_WL 0 0.0748187f
c_342 R1_WL 0 0.082332f
c_371 R3_WL 0 0.0873203f
c_401 R5_WL 0 0.0812971f
c_432 R4_WL 0 0.065704f
c_453 R5_BTLB 0 0.0258078f
c_473 R4_BTLB 0 0.0191587f
c_491 R3_BTLB 0 0.0226316f
c_511 R2_BTL 0 0.0222487f
c_532 R1_BTL 0 0.0214901f
c_550 R3_BTL 0 0.0220319f
c_569 R5_BTL 0 0.0243208f
c_590 R4_BTL 0 0.0216896f
c_609 W4_BTL 0 0.0218473f
c_628 W5_BTL 0 0.0247192f
c_646 W3_BTL 0 0.0208214f
c_663 W1_BTL 0 0.0254001f
c_679 W2_BTL 0 0.0457277f
c_699 qbar_new 0 0.0502936f
c_726 qbar 0 0.17794f
c_756 GND! 0 0.135692f
c_782 VDD! 0 0.116938f
c_801 qnew 0 0.0518334f
c_828 q 0 0.177718f
*
.include "5r5w.pex.netlist.5R5W.pxi"
*
.ends
*
*
