* File: 4r2w_new.pex.netlist
* Created: Sun Oct 25 19:32:01 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt bitcell_4r2w  R1_WL R2_WL R3_WL R4_WL
+ W1_WL W2_WL
+ R1_BTL R1_BTLB R2_BTL R2_BTLB R3_BTL R3_BTLB R4_BTL R4_BTLB
+ W1_BTL W1_BTLB W2_BTL W2_BTLB

* 
MM3 VDD! q qbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 q qbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM51 R4_BTLB R4_WL net90 GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM47 R1_BTLB R1_WL net90 GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM49 R3_BTLB R3_WL qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM41 qbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM48 R2_BTLB R2_WL qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM42 qbar W2_WL W2_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM94 net90 qbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM95 GND! q net105 GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM0 GND! q qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 q qbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM78 R1_BTL R1_WL net105 GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM80 R4_BTL R4_WL net105 GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM40 W1_BTL W1_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM81 R3_BTL R3_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM39 W2_BTL W2_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM79 R2_BTL R2_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
c_13 R4_BTLB 0 0.0403714f
c_34 R4_WL 0 0.0788857f
c_48 R3_BTLB 0 0.0191806f
c_64 R2_BTLB 0 0.0202702f
c_86 R3_WL 0 0.0637533f
c_105 R2_WL 0 0.0990599f
c_125 R1_WL 0 0.0699728f
c_149 W1_WL 0 0.0767329f
c_167 W2_WL 0 0.0632427f
c_182 R1_BTLB 0 0.019113f
c_199 W1_BTLB 0 0.0187655f
c_215 W2_BTLB 0 0.0184775f
c_230 R1_BTL 0 0.0186971f
c_245 W2_BTL 0 0.0175041f
c_262 W1_BTL 0 0.0200724f
c_276 R4_BTL 0 0.0210725f
c_288 R3_BTL 0 0.0407985f
c_304 R2_BTL 0 0.0199084f
c_316 net90 0 0.0253546f
c_333 qbar 0 0.116376f
c_355 GND! 0 0.0855046f
c_375 VDD! 0 0.073848f
c_387 net105 0 0.0221537f
c_406 q 0 0.112549f
*
.include "4r2w_new.pex.netlist.4R2W_NEW.pxi"
*
.ends
*
*
