* File: 2r1w_new.pex.netlist
* Created: Sun Oct 25 19:26:50 2009
* Program "Calibre xRC"
* Version "v2007.3_36.25"
* 
.subckt bitcell_2r1w  R1_WL R2_WL W1_WL
+ R1_BTL R1_BTLB R2_BTL R2_BTLB W1_BTL W1_BTLB
* 
MM0 GND! q qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15
+ PD=4.6e-07 PS=3.9e-07
MM1 q qbar GND! GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14
+ PD=3.9e-07 PS=4.6e-07
MM3 VDD! q qbar VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
MM2 q qbar VDD! VDD! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
MM41 qbar W1_WL W1_BTLB GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM47 R1_BTLB R1_WL qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM48 R2_BTLB R2_WL qbar GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM40 W1_BTL W1_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM78 R1_BTL R1_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
MM79 R2_BTL R2_WL q GND! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
c_10 R1_BTLB 0 0.0271556f
c_21 R2_BTLB 0 0.0271529f
c_33 W1_WL 0 0.0912803f
c_46 R1_WL 0 0.0832923f
c_55 W1_BTLB 0 0.0338891f
c_67 R2_WL 0 0.0961136f
c_76 W1_BTL 0 0.0414779f
c_87 R1_BTL 0 0.0218744f
c_97 R2_BTL 0 0.0200646f
c_109 qbar 0 0.0864049f
c_122 GND! 0 0.0722726f
c_135 VDD! 0 0.0704239f
c_147 q 0 0.088658f
*
.include "2r1w_new.pex.netlist.2R1W_NEW.pxi"
*
.ends
*
*
